`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:      Sungyoon Jung
// Create Date:   2024
// Module Name:   tb_four_bit_adder_struc.v
// Target Module: four_bit_adder_struc.v
//
// Description:   
//    Testbench for verifying the four bit adder.
//
// Test Strategy:
//   Apply random input to verify the four bit adder.
//////////////////////////////////////////////////////////////////////////////////

module tb_four_bit_adder_behav();

  reg
